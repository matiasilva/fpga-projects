module lcd_st7789v3 (
   input  clk,
   output lcd_rst,
   output lcd_rs,
   output lcd_sd,
   output lcd_scl,
   output lcd_cs
);



endmodule
