`define  MADCTL_CMD 8'h36
`define  COLMOD_CMD 8'h3A
`define PORCTRL_CMD 8'hB2
`define   GCTRL_CMD 8'hB7
`define   VCOMS_CMD 8'hBB
`define LCMCTRL_CMD 8'hC0
`define FRCTRL2_CMD 8'hC6
`define   INVON_CMD 8'h21
`define  DISPON_CMD 8'h29
`define   CASET_CMD 8'h2A
`define   RASET_CMD 8'h2B
`define   RAMWR_CMD 8'h2C

